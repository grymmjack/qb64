�P   ˀ� ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                <x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                  0 �   `     �   0 �   `     �   0 �   `     �   0 �  a_  �������������������?�������������������?�������������������?����������������                                                                        A_                                                                           A_     p �   `     �   0 �   `     �   0 �   `     �   0 �  aD  �������������������?�������������������?�������������������?����������������   @                                                                    AD      @                                                                    AD     p �   `     �   0 �   `     �   0 �   `     �   0 �  bD  �������������������?�������������������?�������������������?����������������   @                                                                    "D      @                                                                    "D    
�}���  `     �   0 �   `     �   0 �   `     �   0 �  tD  �������������������?�������������������?�������������������?����������������  
�m�r�                                                                 D     
�m�r�                                                                 D    )yS�)  `     �   0 �   `     �   0 �   `     �   0 �  hD  ��������������������?�������������������?�������������������?����������������  )IR�)                                                                 D     )IR�)                                                                 D    
$y�$  `     �   0 �   `     �   0 �   `     �   0 �  tD  ��������������������?�������������������?�������������������?����������������  
$I�$                                                                 D     
$I�$                                                                 D      0     `     �   0 �   `     �   0 �   `     �   0 �   @   ���݆��u������������?�������������������?�������������������?�������������                                                                                  
"I�"                                                                 "D      0     `     �   0 �   `     �   0 �   `     �   0 �       ���ֆˬu������������?�������������������?�������������������?�������������                                                                                  
)I4R�)                                                                 AD       �   `     �   0 �   `     �   0 �   `     �   0 �       �����,t������������?�������������������?�������������������?����������������                                                                                  
&(ӊr&                                                                 AD      0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                   0 �   `     �   0 �   `     �   0 �   `     �   0 �   `   �������������������?�������������������?�������������������?����������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                <x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x��Ǐ<x�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç8p�Ç                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       >      <   qς �                                          �����                                                                                                                                                                                                                                                              B   "�(   �                                        (��                                                                                                                                                                                                                                                             @   �(                                             (��                                                                                                                                                                                                                                                        �9$�p @sĴ���/Ă'<z*�                                    9��A(��rb]�9�p                                                                                                                                                                                                                                                <�E$� @�$�P�(�$�Ȣ"�+                                     E$�/�t��RQ(�"                                                                                                                                                                                                               @                                 �}T��0@�$�P� �$�(� ��*                      @              }$�(���BRQ=(" x                                               @                                                                                                                                                                                               �AU� @�$�P� �$�(� ��*                                    A%(��n"RQE(2 �                                                                                                                                                                                                                                              �D�� B�#%P �(�#(���j                                     E%(��2��QE(�"�                                                                                                                                                                                                                                                �8��p <s�$�H>q���<y�                                     9$�A���� a^<��x                                                                                                                                                                                        �                                                                          �                                              �                              �                                                                                                                                                                                                                             �          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             @                                                                               @                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         @                                                                               @                                                                               @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �                                                                               �                                                                               �                                                                                                                                                                                                             �                                                                               �                                                                               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �                                             �                                 �                                             �                                 �                                             �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                                             @                                                                             @                                                                                                                                                                                                                     ��                       @                                                     ��                       @                                                                                                                                                                                                           @         ��                       @                                           @         ��                       @                                                                                                                                                                                                           @         ��                       @                                           @         ��                       @                                                                                                                                                                                                           @         ��                       @                                           @         ��                       @                                                                                                                                                                                                           @         ��                     ����                                         @         ��                     ����                                                                                                                                                                                                         @         ��                     ����                                         @         ��                     ����                                                                                                                                                                                                         @         ��                     ?����                                         @         ��                     ?����                                                                                                                                                                ���������                               @         ��                     �������������                               @         ��                     ����                                                                                                                                                                ���������                               @         ��                     ��������������                               @         ��                     �����                                                                                                                                                                ���������                      |         @         ��                    ��������������                      |         @         ��                    �����                                                                                                                                                                ���������                      |         @         ��                    ��������������                      |         @         ��                    �����                                                                                                                                                                ���������                      |         @        ��                    ��������������                      |         @        ��                    �����                                                                                                                                                                ���������                      �         @        ��                    ��������������                      �         @        ��                    �����                                                                                                                                                                ���������                      �      �������     ��                    ��������������                      �      �������     ��                    �����                                                                                                                                                                ���������                      �      �������     ��                    ?��������������                      �      �������     ��                    ?�����                                                                                                                                                                ����������                    �      �������     ��                    ���������������                    �      �������     ��                    �����                                                                                                                                                                ����������                    �      �������     ��                    ����������������                    �      �������     ��                    ������                                                                                                                                                                ����������                    �     �������     ��                   ����������������                    �     �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ����������������                    ��    �������     ��                   ������                                                                                                                                                                ����������                    ��    �������     ��                   ?����������������                    ��    �������     ��                   ?������                                                                                                                                                                �����������                   ��    �������     ��                   �����������������                   ��    �������     ��                   ������                                                                                                                                                                �����������                   ��    �������     ��                   ������������������                   ��    �������     ��                   �������                                                                                                                                                                �����������                   ��    �������     ��                  ������������������                   ��    �������     ��                  �������                                                                                                                                                                �����������                   ��    �������     ��                  ������������������                   ��    �������     ��                  �������                                                                                                                                                                �����������                  ��    �������     ��                  ������������������                  ��    �������     ��                  �������                                                                                                                                                                �����������                  ��    �������     ��                  ������������������                  ��    �������     ��                  �������                                                                                                                                                                �����������                  ��    �������     ?��                  ������������������                  ��    �������     ?��                  �������                                                                                                                                                                �����������                  ��    �������     ?��                  ������������������                  ��    �������     ?��                  �������                                                                                                                                                                ������������                  ��    �������     ?��                  �������������������                  ��    �������     ?��                  �������                                                                                                                                                                ������������                  ��    �������     ?��                  �������������������                  ��    �������     ?��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                ������������                  ��    �������     ��                  �������������������                  ��    �������     ��                  �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            