�P  (#� G �������������������������������������������������������������������������������������������������������������������������                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             ����������������������������� ����������������������������� �                           ������������������������������ �                            �                            �                           ��                            ����������������������������� ����������������������������� �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �     >  �        ��|     ������������������������������ �                           
 �                           
 �       �         �B     ������������������������������ �                           
 �                           
 �       �         �B     ������������������������������ �                           
 �                           
 �     p<�Hy��g���B     ������������������������������ �                           
 �                           
 �     �"�H�+ H� �|     ������������������������������ �                           
 �                           
 �     �"�H�� O���QB     ������������������������������ �                           
 �                           
 �     �"�H"�* H@�1B     ������������������������������ �                           
 �                           
 �     �"�0"�* H� �1B     ������������������������������ �                           
 �                           
 �     p<� y�$G��B     ������������������������������ �                           
 �                           
 �                        ������������������������������ �                           
 �                           
 �         � �              ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �     |        @   ���    ������������������������������ �                           
 �                           
 �     B        @   �     ������������������������������ �                           
 �                           
 �     B        @  "     ������������������������������ �                           
 �                           
 �     B�1����0H�A�
"     ������������������������������ �                           
 �                           
 �     |�J@IS(�QA""     ������������������������������ �                           
 �                           
 �     @�! �IR/�a�A"
"     ������������������������������ �                           
 �                           
 �     @��IR( QA""     ������������������������������ �                           
 �                           
 �     @�JAFR(�I�" �     ������������������������������ �                           
 �                           
 �     @�1��D�' D� ���     ������������������������������ �                           
 �                           
 �                         ������������������������������ �                           
 �                           
 �                         ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ������������������������������ �                           
 �                           
 �                           ��                            ����������������������������� ����������������������������� �                           ������������������������������ �                            �                            �                           ��                             ����������������������������� ����������������������������� �                           ��                             �                             �                             �������������������������������                             �                             �                             �������������������������������                             �                             �                             ������������������������������                              ������������������������������                              ��������������������������������U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                  