�P  �>  P -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����                               �����                               �����             �����             �����    �����    �����                       �����    �����             �����    �����    �����                       �����    �����             �����    �����    �����                       �����    �����             �����    �����    �����                       �����    �����             �����       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P - ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    �����    ���       �@��׿�       �@��׿�       �@��׿�       �@��׿�       ����� �       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�       �@��׿�  P ���������                    ���������                              ���������                              ���������                              ���������                              ���������          ������������������          ������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������p  � p p  � p                     p  � p p  � p           p  � p                               x  � x                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x 0    0 0    0 0    0 H  � H                               x  � x                               x  � x p  � p p  � p           p  � p p  � p p  � p                     p  � p p  � p           p  � p p �����p �����   �����    ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ������������U  UW����U  UW�             ����� ���U  UW����U  UW�          ���������   UUUUP                     ���������                              ���������          ������������������          ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������������������������                    ������������������          ���������?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����������               >        �  ?����������  ?����������               ?����������  ?����������  ?����