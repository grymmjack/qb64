�P   ˀ�                                                                                                                                                                 ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                       ��                      �������������������������������������������������������� ?������������������������������������������������������������������������������������������������������                                                                                                                                       ��                      �������������������������������������������������������� ?������������������������������������������������������������������������������������������������������                                                                                                                                       ��                      �������������������������������������������������������� ?������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                       ?��                      �������������������������������������������������������� ������������������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                                                                    ������������               �����������������������������������������������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������                          ������������               ��        �����          ���������������������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������                          ������������               ��        �����          ���������������������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������         �                ������������               ��        �����          ���������?�����������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������         �                ������������               ��        �����          ���������?�����������������           �����������������������������������������������������������������������������������������������                                                                                 ?��������     �����������         �                ������������               ��        �����          ���������?�����������������           �����������������������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                                                 ?������������ �����������         �                ������������  ��������������           �          ���������?�����������������           ���           ?��������������������������������������������������������������������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ��������������������������                         ��               ����������                          ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ���������������         ������ ������������������                         ��               ����������       ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ������������������������������� ������������������                         ��                                ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ������������������������������� ������������������                         ��                                ��                 ?����������������������������������������������������������� ������������������                                                            ��                  �������������������������� ������������������������������� ������������������                         ��                                ��                 ?����������������������������������������������������������� ������������������                                                                                �������������������������� ����������������������������������������������������                         ��                                                   ?��������������������������������������������������������������������������������                                                                                �������������������������� ����������������������������������������������������                         ��                                                   ?��������������������������������������������������������������������������������                                                                                �������������������������� ����������������������������������������������������                         ��                                                    ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������                                                                                ��������������������������������������������������������������������������������          ��                                                                    �������������������������������������������������������������������������������                                                                                ���������� �������������������������������������������������������������������          ��                                                                    �������������������������������������������������������������������������������                                                                                ���������� �������������������������������������������������������������������          ��                                                                    ������������������������������������������������������ �����������������������                                                                                ���������� ������������������������������������������ �����������������������          ��                                                                    ������������������������������������������������������ �����������������������                                                                                ���������� ������������������������������������������ �����������������������          ��                                                                    ������������������������������������������������������ �����������������������                                                                                ���������� ������������������������������������������ �����������������������          ��                                                                    ������������������������������������������������������ �����������������������                                                                                ���������� ������������������������������������������ �����������������������          ��                                                                    ������������������������������������������������������ �����������������������                                                                                ���������� ������������������������������������������ �����������������������          ��                                                                    ������������������������������������������������������ �����������������������                                                                                ���������� ������������������������������������������ �����������������������          ��               �������������������������                           ������������������������������������������������������ �����������������������                           �������������������������                           ���������� ������������������������������������������ �����������������������          ��               ?�������������������������                           ���������� ������������������������������������������ �����������������������          ��               ?�������������������������                           ���������� ���������������                        �� �����������������������          ��               �������������������������                           ���������� ������������������������������������������ �����������������������          ��               �������������������������                           ���������� ���������������                        �� �����������������������          ��               ��������������������������                           ���������� ���������������?�������������������������� �����������������������          ��               �?������������������������                           ���������� ����������������                      �� �����������������������          ��              ��������������������������                           ���������� ����������������������������������������� �����������������������          ��              �������������������������~                           ���������� ��������������                        ��� �����������������������                          ��                      �                           ������������������������������������������������������� �����������������������                           ��������������������������                           ���������������������������                      @A�� �����������������������                          ��         ���         ��                           �����������������������������                     ��� �����������������������                           ��                     �                           ��������������������������� �����������������������!�� �����������������������                          ��������������������������                           �������������������������������������������������������������������������������                           �������������������������                           ���������������������������          @            �!���������������������������                          �������������������������                           ��������������������������������������������������������������������������������                           ��������������������������                           ���������������������������           @             ���������������������������                          �������������������������                           ��������������������������������������������������������������������������������                           ��������������������������                           ���������������������������           @             ���������������������������                          ��         8           �                           ��������������������������������������������������������������������������������                           ������������  �����������                           ���������������������������           @             ���������������������������                          ��         ;���         ?�                           �����������������������������         <  >         ����������������������������                           ��         8           �                           ��������������������������� ����������  !�������������������������������������                          �������������������������|                           ���������������������������������������  ?��������������������������������������                           ������������  �����������                           ���������������������������           @             ���������������������������                          �?������������������������                           ���������������������������������������  ?��������������������������������������                           ������������  �����������                           ���������������������������           @             ���������������������������              ��������������������������������������������������               ���������������            ������������  ?�����������           ���������������                           ������������  �����������                          ���������������������������           @             ���������������������������              �������������          ;���          ?������������               ���������������������������������������  ?��������������������������������������              ������������������������  �����������������������               ���������������                       @                          ���������������              �������������          ;���          ?������������               ����������������������������          <  >          ?���������������������������              �������������          8            ?�������������              ���������������            �����������  !�����������            ���������������������       ���������������������������������������������������       ������      ��������������������������������  ?�������������������������������                   ������������������������  �����������������������             ���������������|                      @                        �?���������������������       ���������������������������������������������������       ?���������������������}�����������������������  ?���������������������������������������������       }�����������������������  ������������������������       ?������      ���������                      @                        ��������      �������       ���������������������������������������������������       ���������������������������������������������  ?���������������������������������������������       ������������������������  ������������������������       ������      ��������                      @                        ��������      �������       ��                     ;���                     ��       ���������������������������������������������  ?���������������������������������������������       �����������������������  ������������������������       �������       �������� �                     @                        ��������      �������       ��                     ;���                     ��      �����������������������                      <  >                     ������������������������      �                      8                       ��       �������       ������� �����������������������  !�����������������������������       �������       ��������������������������������������������������      ����������������������������������������������  ?����������������������������������������������      ������������������������  ������������������������       �������       �������                       @                          �������       �������       ��������������������������������������������������      ����������������������������������������������  ?����������������������������������������������      ������������������������  ������������������������       �������       �������                       @                          �������       �������       ����������������  �����������  ?�����������������      ����������������������������������������������  ?����������������������������������������������      ������������������������  ������������������������       �������       �������                       @                          �������       �            ����������������     ;���   0  �����������������      �     ���������������������������������������  ?����������������������������������������������      �����������������  ����  ����  ?�����������������       �������       �������                 ���   @      ���                �������       �            |���������������     ;���   0  �����������������      �     ��������������������������������   <  >   ?��������������������������������������      ����������������     8     8  ?�����������������       ������   ���������               �������  !�������              |��������   ���   ?�       �����������������  �����������  ����������������      ��   ���   ���������������������������������  ?���������������������������������   ���   ��      �����������������  ����  ����  ?�����������������       ��   �       �������                 ���   @      ���                �������      ��   ?����������������{����{����  ����  ����  ����{����{����������������   ���   ��      �������{����{�������������������������{����{�������      ��   ���   ��      �������{����{����  ����  ����  ?����{����{�������      ��   �       �������   !B�!B�!B ���   G���   ��� B�!B�!B   �������      ��   ?����������������{����{���������������8�����{����{����������������   ���   ����������������{����{������������������������{����{����������������   ���   ����������������{����{���������������8�?����{����{����������������   �                  !B�!B�!B ���   @      ��� B�!B�!B                 �     �������� �����{����{�����   ?���   0E����{����{��������������    ��   ����������������{����{�����]������������������{����{����������������   ���   ����������������{����{����������������E?����{����{����������������   �                  !B�!B�!B ���   @      ��� B�!B�!B                 �     �������� �����{����{�����   ?���   0E����{����{��������������    �    �������� �����{����{�����]�   ?���   ?������{����{��������������    �    �������� �����{����{�����   ?���   8E?����{����{��������������    �   ?�        �� !B�!B�!B �������  ������� B�!B�!B �        �   ���   ?��������������������������������������E��������������������������   ���   ���������������������������]����������������������������������������   ���   ��������������������������������������E?��������������������������   �                                ���   @      ���                              ��   ?������������             �����  ����E�            ������������   ���   ���������������������������]����������������������������������������   ���   �������������������������������  ����E?��������������������������   �                                ���   ���   ���                              ��   ?������������             ������������E�            ������������   ���   ���������������������������]����������������������������������������   ���   ������������             ������������E?�            ������������   �                 �����������������          ����������������                �               ����������������          0E���������������              ��   ������������             �]���������������            ������������   ���   ������������             ������������E?�            ������������   �                 �����������������          ����������������                �               ����������������          0E���������������              �              ����������������]�          ?�����������������              �              ����������������          8E?���������������              �   ?�����������               �����������������              �����������   ���   ?�������������������������������������8���������������������������   ���   ��������������������������������������������������������������������   ���   �������������������������������������8�?��������������������������   �                                ���          ���                              ��   ?����������������{����{����  �����������  ����{����{����������������   ���   ����������������{����{�������������������������{����{����������������   ���   ����������������{����{����  �����������  ?����{����{����������������   �                  !B�!B�!B ���          ��� B�!B�!B                 ��   ?����������������{����{����  �����������  ����{����{����������������   ���   ����������������{����{�������������������������{����{����������������   ���   ����������������{����{����  �����������  ?����{����{����������������   �                  !B�!B�!B ���          ��� B�!B�!B                 �               �����{����{����            0  ����{����{�����              ��   ����������������{����{�������������������������{����{����������������   ���   ����������������{����{����  �����������  ?����{����{����������������   �                  !B�!B�!B ���          ��� B�!B�!B                 �               �����{����{����            0  ����{����{�����              �              �����{����{�������          ?�������{����{�����              �              �����{����{����            8  ?����{����{�����              �   ?����������� !B�!B�!B ����������������� B�!B�!B �����������   ���   ?���������������������������������������������������������������������   ���   ��������������������������  �����������  ?��������������������������   ���   ��������������������������  �����������  ?��������������������������   �                                ���          ���                              ��   ?���������������������������������������������������������������������   ���   �������������������������������      �������������������������������   ���   �������������������������������      �������������������������������   �                                    ?�������                                   ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                                                                               ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                       |                                �                     ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                       @                                �                     ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                       @             !<�x           � �                     ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                       @�q�          1B�D           ��                     ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                       y�           1BD�B           L��                     ��   ?���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   ���   ���������������������������������������������������������������������   �                       A��          )BD�B           H��                     ��   ?���������������������������������������������������������������������   ���   �������������������}�����������������������������7]_�����������������   ���   �������������������}�����������������������������7]_�����������������   �                       A�           )BD�B           Ȣ�                     ��   ?���   �������������������������������������������������������   ����   ���   �������������������u�����������ڽ�WZ��������������]]�����������������   ���   �������������������u�����������ڽ�WZ��������������]]�����������������   �                       A�           %B��B           (��                     ��   ?���������������������������������������������������������������������   ���   �������������������?����������ܽ�W\��������������ac�����������������   ���   �������������������?����������ܽ�W\��������������ac�����������������   �                      @�q�          #B��B           (��                    ��   ?���   �������������������������������������������������������  ����   ���   �������������������������������ܽ��\���������������������������������   ���   ���   ������������������������ܽ��\��������������������������  ����   �         ����                        #B�D                       ���        ��   ?��������������������������������������������������������������������   ���   �����������������������������������^���������������������������������   ���   ����������������������������������^���������������������������������   �         �  (                        !<�x             <                    ���������������������������������������������������������������������������������   ���������������������������������������������������������������������   ���   ��������������������������������������������������������������������   � ����   �  (                                                           ���� ���������   �������������������������������������������������������  ������������������   �������������������������������������������������������  ������������������   �������������������������������������������������������  ���������         ����                                                      ���         ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                              ���������   ������������������������      ������������������������   ������������������   �������������������������������������������������������   ������������������   �������������������������������������������������������   ���������        ����                                                      ?���         �������������������������������������      ���������������������������������������������������������������������������������������������������������������������������������������������������������      ������������������������������������                                    ?�������                                    ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            