�P   N � ���������������������������������������������������������������������������������������������������������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �?������������������������������?����������������������������� ��                            ������������������������������� �                             �                              ��                            ��                             �/������������������������������/����������������������������� ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                        ����(�(                        ����( ��                        ���������������������������������� �(                        ����(�(                        ����( ��                        �������������������������������?�� �( �9��O>�Bp              ����(�( �9��O>�Bp              ����( �� �9��O>�Bp              ��?���������������������������� �� �( �DD(P��b�              ����(�( �DD(P��b�              ����( �� �DD(P��b�              � ���������������������������� �� �( �@D(P�b�              ����(�( �@D(P�b�              ����( �� �@D(P�b�              � ���������������������������� �� �( �@D(P�R�              ����(�( �@D(P�R�              ����( �� �@D(P�R�              � ���������������������������� �� �(                        �� (�(                        �� ( �� �8G�P�Rp              � ���������������������������� �� �(                        �� (�(                        �� ( �� �D(P�J              � ���������������������������� �� �(                        �� (�(                        �� ( �� �D(P�F              � ���������������������������� �� �(                        �� (�(                        �� ( �� �DD(P��F�              � �����������������������������?�� �(                          � (�(                          � ( �� �8D'��Bp              ��?������������������������������� �(                          � (�(                          � ( ��                        ���������������������������������� �(                            (�(                            ( ��                        ����������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( �� �(       @    @         ������������������������������ �(                            (�(                            ( �� �(       @    @ H        ������������������������������� �(                            (�(                            ( �� DH       @    @ H        ������O������c*������m������� �(                            (�(                            ( �� DK�'s��8X�k3�N`    �����]7��_mu��]j��}��[�������� �(                            (�(                            ( �� DL��������eL�RQ@    ����wAw��Xm��]j�����[�������� �(                            (�(                            ( �� *��������<E�H�U_@    ����w_w��Wm}��]j������[�������� �(                            (�(                            ( �� *���"�����DE H�UP@    �����]w��Wsu��]j��}��[�n������ �(                            (�(                            ( �� ��"�����D�EH�H�@    �����cw���w���cj�����\wq������ �(                            (�(                            ( �� ��'�r��<D�(���D    ������������������������������ �(                            (�(                            ( ��          �              ������������������������������� �(                            (�(                            ( ��       0                  ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( ��  }� *         �       ���o��������������������������� �(                            (�(                            ( �� � A 
              @  ���o��������������������������� �(                            (�(                            ( �� � A 
              @  ���)�����U���Lq��g�g��'�Ӈ�� �(                            (�(                            ( �� �8A$���XX�,�9��G,x ���f�����U�]�[�����[����Mw�� �(                            (�(                            ( �� �Dy$���QdeP2�%@�� ���n�����U�A�X ���/�o����]w�� �(                            (�(                            ( �� �|A*����DE�"�=%�G�� ���n�����U�_�[�����w����]w�� �(                            (�(                            ( �� �@A*���DE"�E% H�� ���n�������]�[�����[���]w�� �(                            (�(                            ( �� �DA*��QDEP"�E%H�� �������������\q��o�g����]��� �(                            (�(                            ( �� Q8}�*��DD�"�=$�G�x ������������������������������ �(                            (�(                            ( ��           �            @   ������������������������������� �(                            (�(                            ( ��                           ������������������������������� �(                            (�(                            ( ��                            ����}����_�������������������� �(                            (�(                            ( �� �
�   �       (   @    ����}�������������_���������� �(                            (�(                            ( �� �
�   �      �  @    ����}������������������������ �(                            (�(                            ( �� �
�   �         @    ���N=|8�8�T���8Ӎ8���6�4������ �(                            (�(                            ( �� ���'��,r�)��X�   ���5�}�|�WS]�}�M��o�����}������ �(                            (�(                            ( �� �"�(�(��� � � �**,�e   ���t}�}�WW]�}�]��o�����}����� �(                            (�(                            ( �� ��/�(����'�z'�*(�E�   ���u�}���WW]�}�]u�o�����}������ �(                            (�(                            ( �� ��((����(��(�*
(�E    ���u�}�}�WW]�}�]u�o�U���}������ �(                            (�(                            ( �� �"�(�(����(��(��)(�E   ���v=|8���Wa�|8]��k��7~7~����� �(                            (�(                            ( �� ��''���Ǣz'�)ȁȁD�   ������������������������������� �(                            (�(                            ( ��                          ������������������������������� �(                            (�(                            ( ��         <                  ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��              @@ ����������������������߷������� �(                            (�(                            ( ��            H   @ ����������������������߷������� �(                            (�(                            ( �� (           H   @ ����������Ӈ�1����
�ϔ��4���� �(                            (�(                            ( �� (���e<�,x�<�8�0k
�N@ �������j���Mw�~�������_�]�վ��� �(                            (�(                            ( �� D�* �E ��"�D	�L�*A@ ����������]w�p�������߷A�հ��� �(                            (�(                            ( �� D�+�EE���"�D	= H�
*O@ �������ں��]w�n������߷_�ծ��� �(                            (�(                            ( �� |�* %E��"�D	E H�
*Q@ �������j���]w�n������_�]�ծ��� �(                            (�(                            ( �� ��* �E��"�D	E4�H�
*Q@ ����������]��p����,��c�ְ��� �(                            (�(                            ( �� ����e<��x�<�<��(�
)O@ ������������������������������� �(                            (�(                            ( ��                          ������������������������������� �(                            (�(                            ( ��  �         x             ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( ��        �    @     @  ���o��������ۿ���������������� �(                            (�(                            ( �� �       $@          �@  ���o��������ۿ���������������� �(                            (�(                            ( �� �       $@          �@  ���)��T��Ӆ�ۿp�㟳��8��1���� �(                            (�(                            ( �� �g$�,zp$@�g`L�5�,�@  ���f�[S]�Muw۾뮷]o��|�[�M~���� �(                            (�(                            ( �� �H��� ���$AQH��R �(�(��@  ���n�UW]�]u۾�.�A���}�[�]p���� �(                            (�(                            ( �� �H������$A�O�@H�(�H��@  ���n�UW]�]u۾���߻�}�[w]n���� �(                            (�(                            ( �� �H������$AH  D�(����@  ���n�n�]�]uw۾뮷]o��}�Z�]n���� �(                            (�(                            ( �� �H�(����$AQH��R�(���@  �������a�]���p�㟳�}��ݰ���� �(                            (�(                            ( �� QG(��zp#��G`L�'%�"O@  ������������������������������� �(                            (�(                            ( ��                         ������������������������������ �(                            (�(                            ( ��     <  �                 ������������������������������� �(                            (�(                            ( ��                            ����������������W�������������� �(                            (�(                            ( ��          �   @ p    ���o��������������������w����� �(                            (�(                            ( �� �    $      (    ��   ���o������������������������� �(                            (�(                            ( �� �    $      (    ��   ���)��}O�q�e8��V>
c���~3���� �(                            (�(                            ( �� �g$��5���0<�����sNX���   ���f�[}7ٮ���_��Wݾ��u�������� �(                            (�(                            ( �� �H���&QS(�E�"A"�Qd�r(   ���n�U}w۠���_��V���}������� �(                            (�(                            ( �� �H���$_R/�E��>�QD��   ���n�U}wۯ���ߺ�U�~��}�������� �(                            (�(                            ( �� �H���$PR( E� � �QD�
   ���n�n�wۮ���_��Uݾ��u��u����� �(                            (�(                            ( �� �H��$QR(�E�"A"�QD��(   �������w��u���V
㎱�_�;���� �(                            (�(                            ( �� QG�N�' <���qND�q�   ������������������������������ �(                            (�(                            ( ��                     �     ������������������������������� �(                            (�(                            ( ��            x              ������������������������������� �(                            (�(                            ( ��                            ������������������������������ �(                            (�(                            ( ��     A          �     ���o��������������������������� �(                            (�(                            ( �� �       $             ���o��������������������������� �(                            (�(                            ( �� �       $             ���)�������}O�q����c�������� �(                            (�(                            ( �� �89�pO9��5��p$�H�  ���f�����ڮ��7ٮ�}mw�}�����[��� �(                            (�(                            ( �� �DE"�%QE�&Q���$�H"	�  ���n������w۠��m�a��������� �(                            (�(                            ( �� �|E �Q}�$_��*�H"	  ���n���������wۯ��m�]��������� �(                            (�(                            ( �� �@E �	QA�$P"��*�H"	  ���n�����ڮ��wۮ�]mw�������[��� �(                            (�(                            ( �� �DE"�%QE�$Q���"0"	�  ������������w���m����������� �(                            (�(                            ( �� Q89pO9�N�p"�  ������������������������������� �(                            (�(                            ( ��                            ����������������������?�������� �(                            (�(                            ( ��                    �       ������������������������������� �(                            (�(                            ( ��                            �������������������������� ���� �(                            (�(                            ( ��       
              ���o����������o����������� ���� �(                            (�(                            ( �� �       �            ���o����������o����������� ���� �(                            (�(                            ( �� �       �            ���)��Ɯi��5��)�������Li� ���� �(                            (�(                            ( �� �89c�8�r@�89c�8E��     ���f���o����uf�������ۦ� ���� �(                            (�(                            ( �� �D�Y*���D�YE$Y     ���n����.���|�n�������ۮ� ���� �(                            (�(                            ( �� �|=�<
� �|=�<E$Q     ���n��뮻��}n�������ۮ� ���� �(                            (�(                            ( �� �@EQD
���@EQDE$Q     ���n��뮻��u�n�������ۮ� ���� �(                            (�(                            ( �� �DEQD*�@�DEQDM$Q     ��������.�~5�߮��������ln� ���� �(                            (�(                            ( �� Q8=�<��r Q8=�<4��     �������������������������� ���� �(                            (�(                            ( ��                           �������������������������� ���� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ������������������������������� �(                            (�(                            ( ��                            ��                             �/������������������������������/����������������������������� ��                            ������������������������������� �                             �                              ��                            ��                               �?������������������������������?����������������������������� ��                            ��                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ���������������������������������                               �                              �                               ��������������������������������                                ��������������������������������                                ��������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            